class jk_transaction;
    rand logic J, K;  // Randomize values for J and K

    // Constructor
    function new();
        J = 0;
        K = 0;
    endfunction
endclass
